*$
* INA849
*****************************************************************************
* (C) Copyright 2022 Texas Instruments Incorporated. All rights reserved.
*****************************************************************************
** This model is designed as an aid for customers of Texas Instruments.
** TI and its licensors and suppliers make no warranties, either expressed
** or implied, with respect to this model, including the warranties of
** merchantability or fitness for a particular purpose.  The model is
** provided solely on an "as is" basis.  The entire risk as to its quality
** and performance is with the customer
*****************************************************************************
*
* This model is subject to change without notice. Texas Instruments
* Incorporated is not responsible for updating this model.
*
*****************************************************************************
*
** Released by: Online Design Tools, Texas Instruments Inc.
* Part: INA849
* Date: 18JUL2022
* Model Type: Generic (suitable for all analysis types)
* EVM Order Number: NA
* EVM Users Guide:  NA
* Datasheet: SBOS945B – NOVEMBER 2020 – REVISED APRIL 2021
* Created with Green-Williams-Lis Op Amp Macro-model Architecture
*
* Model Version: Final 1.1
*
*****************************************************************************
*
*
* Updates:
*
* Final 1.1
* 1. Updated PSpice Symbol.
* 2. Added .ENDS name as INA849.
* 3. Moved R_NOISELESS .model inside INA849 Subckt.
*
* Final 1.0
* Release to Web.
* INA849 - Rev. A
* Created by Srivatsan Sathyamoorthy; 2020-12-08
* Created with Green-Williams-Lis Current Sense Amp Macro-model Architecture
* Copyright 2020 by Texas Instruments Corporation
*
*****************************************************************************
* MACRO-MODEL SIMULATED PARAMETERS:
*****************************************************************************
* AC PARAMETERS
*****************************************************************************
* CLOSED-LOOP OUTPUT IMPEDANCE VS. FREQUENCY (Zout vs. Freq.)
* CLOSED-LOOP GAIN AND PHASE VS. FREQUENCY  WITH RL, CL EFFECTS (Acl vs. Freq.)
* COMMON-MODE REJECTION RATIO VS. FREQUENCY (CMRR vs. Freq.)
* POWER SUPPLY REJECTION RATIO VS. FREQUENCY (PSRR vs. Freq.)
* INPUT VOLTAGE NOISE DENSITY VS. FREQUENCY (en vs. Freq.)
*****************************************************************************
* DC PARAMETERS
*****************************************************************************
* INPUT COMMON-MODE VOLTAGE RANGE (Vcm)
* GAIN ERROR (Eg)
* INPUT BIAS CURRENT VS. INPUT COMMON-MODE VOLTAGE (Ib vs. Vcm)
* INPUT OFFSET VOLTAGE VS. TEMPERATURE (Vos vs. Temp)
* OUTPUT VOLTAGE SWING vs. OUTPUT CURRENT (Vout vs. Iout)
* SHORT-CIRCUIT OUTPUT CURRENT (Isc)
* QUIESCENT CURRENT (Iq)
*****************************************************************************
* TRANSIENT PARAMETERS
*****************************************************************************
* SLEW RATE (SR)
* SETTLING TIME VS. CAPACITIVE LOAD (ts)
*****************************************************************************
* CONNECTIONS:  NON-INVERTING INPUT
*               |   INVERTING INPUT
*               |   |   POSITIVE POWER SUPPLY
*               |   |   |   NEGATIVE POWER SUPPLY
*               |   |   |   |   OUTPUT
*               |   |   |   |   |    REFERENCE
*               |   |   |   |   |    |   GAIN SET 1
*               |   |   |   |   |    |   |   GAIN SET 2
*               |   |   |   |   |    |   |   |
.SUBCKT INA849  IN+ IN- VCC VEE OUT REF RG+ RG-
*****************************************************************************
C_C13            0 N1602505  1F
C_C14            0 N1602365  10N
C_C15            0 N1602545  1F
C_C16            N1604573 REF  1F
C_C17            N1604535 OUT  11F
C_CCM1           MID INP  1F
C_CCM2           MID INN  1F
C_CIN_CMN        ESDN MID  7P
C_CIN_CMP        MID ESDP  7P
C_C_GS1          NODE1 N969492  2.6P
C_C_GS2          NODE2 N969473  2.6P
E_E_MID          MID 0 N1602365 0 1
G_GM1            N969492 RG- INN RG- 22.02M
G_GM2            N969473 RG+ INP RG+ 22.02M
G_G_VCC_BUFFER   VCC_B 0 VCC 0 -1
G_G_VEE_BUFFER   VEE_B 0 VEE 0 -1
I_IB             N1383401 MID DC 10PADC
I_IOS            N1383384 MID DC 5PADC
I_I_Q            VCC VEE DC 6.2M
I_I_SINK1        RG- VEE_B DC 24UADC
I_I_SINK2        RG+ VEE_B DC 24UADC
R_RCM1           MID N1385067 R_NOISELESS 1T
R_RCM2           N1385271 MID R_NOISELESS 1T
R_RCM3           N1385582 MID R_NOISELESS 1
R_RCM4           N1385582 INP R_NOISELESS 1M
R_RCM5           MID N1386246 R_NOISELESS 1T
R_RCM6           N1386314 INN R_NOISELESS 1M
R_RCM7           N1386314 MID R_NOISELESS 1
R_RCM8           N1386438 MID R_NOISELESS 1T
R_RF1            RG- NODE1  3K
R_RF2            RG+ NODE2  3K
R_RFN            N1604535 OUT  5.0000316K
R_RFP            N1604573 REF  5K
R_RIN11          ESDP IN+ R_NOISELESS 10M
R_RIN12          ESDN IN- R_NOISELESS 10M
R_RIN13          N1384907 N1384032 R_NOISELESS 10M
R_RIN14          N1386364 N1383384 R_NOISELESS 10M
R_RIN_CMN        MID ESDN R_NOISELESS 1T
R_RIN_CMP        ESDP MID R_NOISELESS 1T
R_RIN_IN         NODE1 N1604535  5K
R_RIN_NIN        NODE2 N1604573  5K
R_R_GS1          N969492 VCC_B  41.67K
R_R_GS2          N969473 VCC_B  41.67K
R_R_MID1         VCC_B 0 R_NOISELESS 1
R_R_MID2         VEE_B 0 R_NOISELESS 1
R_R_MID3         VCC_B N1602505 R_NOISELESS 1M
R_R_MID4         N1602545 VEE_B R_NOISELESS 1M
R_R_MID5         N1602505 N1602365 R_NOISELESS 1MEG
R_R_MID6         N1602365 N1602545 R_NOISELESS 1MEG
R_R_MID7         N1602365 0 R_NOISELESS 1T
V_VB             VCC_B N969449 1VDC
V_VCM_MAX        N1385067 VCC_B -2.5VDC
V_VCM_MAX1       N1386246 VCC_B -2.5VDC
V_VCM_MIN        N1385271 VEE_B 2.5VDC
V_VCM_MIN1       N1386438 VEE_B 2.5VDC
X_INA849_INAMP0  N969449 N969492 MID VCC VEE NODE1 INA849_INAMP
X_INA849_INAMP1  N969449 N969473 MID VCC VEE NODE2 INA849_INAMP
X_INA849_OUTAMP  N1604573 N1604535 VCC VCC_B VEE VEE_B MID OUT INA849_OUTAMP
X_U1             ESDP N1383401 VNSE1_INA849 PARAMS:  FLW=100M NLF=9 NVR=0.7
X_U10            N1384907 MID N1385582 MID N1385067 N1385271 VCM_CLAMP_INA849 PARAMS:
+  GAIN=1
X_U11            N1386364 MID N1386314 MID N1386246 N1386438 VCM_CLAMP_INA849 PARAMS:
+  GAIN=1
X_U12            RG- VCC VEE ESD_OUT_INA849
X_U13            RG+ VCC VEE ESD_OUT_INA849
X_U14            REF VCC VEE ESD_OUT_INA849
X_U15            OUT VCC VEE ESD_OUT_INA849
X_U16            ESDN N1383384 VNSE1_INA849 PARAMS:  FLW=100M NLF=9 NVR=0.7
X_U3             ESDP VCC VEE ESD_OUT_INA849
X_U4             ESDN VCC VEE ESD_OUT_INA849
X_U7             MID N1383401 FEMT2_INA849 PARAMS: FLWF=0.1 NLFF=17K NVRF=1.06K
X_U8             N1383384 MID FEMT2_INA849 PARAMS: FLWF=0.1 NLFF=17K NVRF=1.06K
X_U9             N1384032 N1383401 VOS_DRIFT_INA849 PARAMS:  DC=10U POL=1 DRIFT=100N
.MODEL R_NOISELESS RES (T_ABS=-273.15)
.ENDS  INA849
*
.SUBCKT ESD_OUT_INA849 OUT VCC VEE
.MODEL ESD_SW VSWITCH(RON=50 ROFF=1E12 VON=500E-3 VOFF=100E-3)
S1 VCC OUT OUT VCC ESD_SW
S2 OUT VEE VEE OUT ESD_SW
.ENDS  ESD_OUT_INA849
*
.SUBCKT FEMT2_INA849  1 2 PARAMS: NLFF = 0.1 FLWF = 0.001 NVRF = 0.1
.PARAM GLFF={PWR(FLWF,0.25)*NLFF/1164}
.PARAM RNVF={1.184*PWR(NVRF,2)}
.MODEL DVNF D KF={PWR(FLWF,0.5)/1E11} IS=1.0E-16
I1 0 7 10E-3
I2 0 8 10E-3
D1 7 0 DVNF
D2 8 0 DVNF
E1 3 6 7 8 {GLFF}
R1 3 0 1E9
R2 3 0 1E9
R3 3 6 1E9
E2 6 4 5 0 10
R4 5 0 {RNVF}
R5 5 0 {RNVF}
R6 3 4 1E9
R7 4 0 1E9
G1 1 2 3 4 1E-6
C1 1 0 1E-15
C2 2 0 1E-15
C3 1 2 1E-15
.ENDS  FEMT2_INA849
*
.SUBCKT VCM_CLAMP_INA849 VIN+ VIN- IOUT- IOUT+ VP+ VP- PARAMS: GAIN=1
G1 IOUT+ IOUT- VALUE={LIMIT(GAIN*V(VIN+,VIN-),V(VP-,VIN-), V(VP+,VIN-))}
.ENDS  VCM_CLAMP_INA849
*
.SUBCKT VNSE1_INA849 1 2 PARAMS: FLW=1 NLF=120 NVR=18
.PARAM GLF={PWR(FLW,0.25)*NLF/1164}
.PARAM RNV={1.184*PWR(NVR,2)}
.MODEL DVN D KF={PWR(FLW,0.5)/1E11} IS=1.0E-16
I1 0 7 10E-3
I2 0 8 10E-3
D1 7 0 DVN
D2 8 0 DVN
E1 3 6 7 8 {GLF}
R1 3 0 1E9
R2 3 0 1E9
R3 3 6 1E9
E2 6 4 5 0 10
R4 5 0 {RNV}
R5 5 0 {RNV}
R6 3 4 1E9
R7 4 0 1E9
E3 1 2 3 4 1
.ENDS  VNSE1_INA849
*
.SUBCKT VOS_DRIFT_INA849 VOS+ VOS- PARAMS: DC=496.4E-6 POL=1 DRIFT=2E-06
E1 VOS+ VOS- VALUE={DC+POL*DRIFT*(TEMP-27)}
.ENDS  VOS_DRIFT_INA849
*$
*
*****************************************************************************
.SUBCKT INA849_OUTAMP OUP_IN+ OUP_IN- VCC VCC_B VEE VEE_B MID OUP_OUT
*****************************************************************************
C_C106          N1661226 MID  1F
C_C107          MID N1661626  1F
C_C108          N1661462 MID  1P
C_C109          MID N1661680  1P
C_C110          N1663763 MID  1P
C_C111          MID N1664091  1P
C_C112          N1663947 MID  1P
C_C113          MID N1664179  1P
C_C114          VCLP MID  1P
C_C115          N1939474 N1939484  418U
C_C116          N1939514 N1939524  324F
C_C117          N1939534 N1939542  31.83F
C_C118          N1939552 N1939562  31.83F
C_C119          N1939572 N1939580  31.83F
C_C120          MID N1940758  2.49P
C_C121          MID N1940790  2.49P
C_C122          MID N1940844  26.98F
C_C123          MID N1940876  26.98F
C_C13           N1939494 N1939504  723N
C_C29           N1428789 N1428799  677F
C_C30           N1428809 N1428819  677F
C_C33           CLAMP MID  900N
C_C34           MID N1428991  13.5F
C_CCM2          MID N995776  1F
C_CIN2_CMN      N953203 MID  1P
C_CIN2_CMP      MID N953165  1P
C_CIN2_DIFF     N953165 N953203  1P
C_CP1           N1389051 N1389061  144.7P
C_CP2           MID N1389297  26.53F
C_CP3           N1388079 N1388089  41.88P
C_CP4           N1388099 N1388109  13.26P
C_CP5           N1388119 N1388129  13.26P
C_CP6           MID N1388615  79.58F
C_CP7           MID N1388629  79.58F
C_C_VIMON       VIMON MID  1P
C_C_VOUTS       VOUT_S MID  1P
E_E2            N1696516 MID CL_CLAMP_OP MID 1
E_E4            N1403176 MID OUP_OUT MID 1
G_G18           N1939722 MID N1939504 MID -114.5
G_G53           VCC_CLP MID N1661226 MID -1M
G_G57           N1394772 N1394706 PSRR+ PSRR- -1M
G_G58           CLAW_CLAMP_OP MID N1428819 MID -1M
G_G59           CL_CLAMP_OP MID CLAW_CLAMP_OP MID -1M
G_G60           N1428789 MID N1428991 MID -6.381
G_G61           N1428809 MID N1428799 MID -6.381
G_G64           VSENSE MID CLAMP MID -1E-3
G_G65           N1428991 MID VSENSE MID -1E-6
G_G66           VEE_CLP MID N1661626 MID -1M
G_G69           N1939474 MID CL_CLAMP_OP OUT_NODE -89
G_G70           N1939494 MID N1939484 MID -1.316K
G_G71           N1939792 MID N1939524 MID -1.63
G_G72           N1939552 MID N1939542 MID -20
G_G73           N1939572 MID N1939562 MID -20
G_G74           N1939746 MID N1939730 MID -1
G_G75           N1939514 MID N1939754 MID -1
G_G76           N1939816 MID N1939800 MID -1
G_G77           N1939534 MID N1939824 MID -1
G_G_PSRNEG      N1388079 MID VEE_B MID -10.53M
G_G_PSRNEG1     N1388099 MID N1388089 MID -1
G_G_PSRNEG2     N1388119 MID N1388109 MID -16.67
G_G_PSRNEG3     N1388139 MID N1388129 MID -16.67
G_G_PSRNEG4     N1388167 MID N1388149 MID -1
G_G_PSRNEG5     PSRR- MID N1388177 MID -1
G_G_PSRPOS      N1389051 MID VCC_B MID -1.818
G_G_PSRPOS1     N1389071 MID N1389061 MID -1
G_G_PSRPOS2     PSRR+ MID N1389081 MID -1
R_R120          N1661302 VCC_B R_NOISELESS 1K
R_R121          VEE_B N1661612 R_NOISELESS 1K
R_R122          N1661226 N1661302 R_NOISELESS 1
R_R123          N1661626 N1661612 R_NOISELESS 1
R_R124          VCC_CLP MID R_NOISELESS 1K
R_R125          MID VEE_CLP R_NOISELESS 1K
R_R126          VCC_CLP MID R_NOISELESS 1T
R_R127          MID VEE_CLP R_NOISELESS 1T
R_R128          N1661466 MID R_NOISELESS 1
R_R129          MID N1661666 R_NOISELESS 1
R_R130          N1661462 N1661466 R_NOISELESS 1
R_R131          N1661680 N1661666 R_NOISELESS 1
R_R142          MID N1664165 R_NOISELESS 1
R_R143          MID N1664265 R_NOISELESS 1G
R_R145          N1394772 N1394706 R_NOISELESS 1K
R_R146          MID CLAW_CLAMP_OP R_NOISELESS 1K
R_R147          MID CL_CLAMP_OP R_NOISELESS 1K
R_R148          N1428799 N1428789 R_NOISELESS 10K
R_R149          N1428819 N1428809 R_NOISELESS 10K
R_R152          MID N1428789 R_NOISELESS 1
R_R153          MID N1428809 R_NOISELESS 1
R_R156          N1428991 MID R_NOISELESS 1E6
R_R157          MID N1428799 R_NOISELESS 1.858K
R_R158          MID N1428819 R_NOISELESS 1.858K
R_R161          MID VSENSE R_NOISELESS 1E3
R_R162          N1663647 MID R_NOISELESS 1T
R_R163          N1663665 MID R_NOISELESS 1G
R_R164          N1663805 MID R_NOISELESS 1
R_R165          N1663951 MID R_NOISELESS 1
R_R166          N1663763 N1663805 R_NOISELESS 1
R_R167          N1663947 N1663951 R_NOISELESS 1
R_R168          N1664091 N1664077 R_NOISELESS 1
R_R169          N1664179 N1664165 R_NOISELESS 1
R_R170          MID N1664077 R_NOISELESS 1
R_R171          MID N1664201 R_NOISELESS 1T
R_R172          N1939730 N1939722 R_NOISELESS 25.56K
R_R173          N1939754 N1939746 R_NOISELESS 25.56K
R_R174          N1939800 N1939792 R_NOISELESS 49K
R_R175          N1939824 N1939816 R_NOISELESS 49K
R_R176          N1939484 N1939474 R_NOISELESS 10K
R_R177          N1939524 N1939514 R_NOISELESS 10K
R_R178          N1939542 N1939534 R_NOISELESS 10K
R_R179          N1939562 N1939552 R_NOISELESS 10K
R_R180          N1939580 N1939572 R_NOISELESS 10K
R_R181          N1940758 N1939730 R_NOISELESS 10K
R_R182          N1940790 N1939754 R_NOISELESS 10K
R_R183          N1940844 N1939800 R_NOISELESS 10K
R_R184          N1940876 N1939824 R_NOISELESS 10K
R_R185          MID N1939722 R_NOISELESS 1
R_R186          MID N1939792 R_NOISELESS 1
R_R187          MID N1939816 R_NOISELESS 1
R_R188          MID N1939534 R_NOISELESS 1
R_R189          MID N1939552 R_NOISELESS 1
R_R190          MID N1939572 R_NOISELESS 1
R_R191          MID N1940296 R_NOISELESS 1
R_R192          MID N1939474 R_NOISELESS 1
R_R193          MID N1939484 R_NOISELESS 7.606
R_R194          MID N1939524 R_NOISELESS 15.81K
R_R195          MID N1939542 R_NOISELESS 526.3
R_R196          MID N1939562 R_NOISELESS 526.3
R_R197          MID N1939580 R_NOISELESS 526.3
R_R198          MID N1939746 R_NOISELESS 1
R_R199          MID N1939514 R_NOISELESS 1
R_R37           MID N1939494 R_NOISELESS 1
R_R44           N1939504 N1939494 R_NOISELESS 10K
R_R45           MID N1939504 R_NOISELESS 88.07
R_R84           N1696516 VCLP R_NOISELESS 100
R_RCM5          MID N1401129 R_NOISELESS 1T
R_RCM6          N1401213 N995776 R_NOISELESS 1M
R_RCM7          N1401213 MID R_NOISELESS 1
R_RCM8          N1401349 MID R_NOISELESS 1T
R_RDUMMY        MID OUT_NODE R_NOISELESS 50K
R_RIN2_CMN      MID N953203 R_NOISELESS 1T
R_RIN2_CMP      N953165 MID R_NOISELESS 1T
R_RIN3          N953165 OUP_IN+ R_NOISELESS 10M
R_RIN4          N953203 OUP_IN- R_NOISELESS 10M
R_RO1           MID N261787 R_NOISELESS 1MEG
R_RO2           MID CLAMP R_NOISELESS 1MEG
R_RP1           N1389061 N1389051 R_NOISELESS 100MEG
R_RP10          N1388129 MID R_NOISELESS 638.3
R_RP11          N1388139 N1388149 R_NOISELESS 90K
R_RP12          N1388149 N1388615 R_NOISELESS 10K
R_RP13          N1388167 N1388177 R_NOISELESS 90K
R_RP14          N1388177 N1388629 R_NOISELESS 10K
R_RP2           N1389061 MID R_NOISELESS 55
R_RP3           N1389071 N1389081 R_NOISELESS 290K
R_RP4           N1389081 N1389297 R_NOISELESS 10K
R_RP5           N1388089 N1388079 R_NOISELESS 100MEG
R_RP6           N1388089 MID R_NOISELESS 9.5K
R_RP7           N1388109 N1388099 R_NOISELESS 10K
R_RP8           N1388109 MID R_NOISELESS 638.3
R_RP9           N1388129 N1388119 R_NOISELESS 10K
R_RSRC          MID N1389051 R_NOISELESS 1
R_RSRC1         MID N1389071 R_NOISELESS 1
R_RSRC2         MID PSRR+ R_NOISELESS 1
R_RSRC3         MID N1388079 R_NOISELESS 1
R_RSRC4         MID N1388099 R_NOISELESS 1
R_RSRC5         MID N1388119 R_NOISELESS 1
R_RSRC6         MID N1388139 R_NOISELESS 1
R_RSRC7         MID N1388167 R_NOISELESS 1
R_RSRC8         MID PSRR- R_NOISELESS 1
R_RX            OUT_NODE N1940296 R_NOISELESS 500K
R_R_VIMON21     MID N989282 R_NOISELESS 1T
R_R_VIMON22     N989282 VIMON R_NOISELESS 100
R_VOUTS1        MID N1403176 R_NOISELESS 1T
R_VOUTS2        VOUT_S N1403176 R_NOISELESS 100
V_VCM_MAX2      N1401129 VCC_B -2VDC
V_VCM_MIN2      N1401349 VEE_B 2VDC
V_V_GRN         N1664265 MID -220VDC
V_V_GRP         N1663665 MID 220VDC
V_V_ISCN        N1664201 MID -34VDC
V_V_ISCP        N1663647 MID 34VDC
X_H_IMON        OUT_NODE OUP_OUT N989282 MID OUTAMP_BLOCK_DC_H_IMON_INA849_OUTAMP
X_U1            N953165 N2052331 VNSE1_INA849_OUTAMP PARAMS:  FLW=150M NLF=524.25 NVR=21
X_U10           N1394772 MID N1401213 MID N1401129 N1401349 VCM_CLAMP_INA849_OUTAMP PARAMS:
+  GAIN=1
X_U11           VIMON MID N1661302 VCC_B CLAWP_INA849_OUTAMP
X_U12           MID VIMON VEE_B N1661612 CLAWN_INA849_OUTAMP
X_U13           VCC_CLP VEE_CLP VOUT_S MID N1661466 N1661666 CLAMP_AMP_LO_INA849_OUTAMP PARAMS:
+   G=25
X_U14           N1661462 N1661680 CLAW_CLAMP_OP MID CLAW_SRC_INA849_OUTAMP PARAMS:  GAIN=1
+  IPOS=500M INEG=-500M
X_U15           N1663647 N1664201 VOUT_S MID N1663805 N1664077 CLAMP_AMP_LO_INA849_OUTAMP
+  PARAMS:  G=25
X_U16           N1663763 N1664091 CL_CLAMP_OP MID CL_SRC_INA849_OUTAMP PARAMS:  GAIN=1 IPOS=1
+  INEG=-1
X_U17           N1663665 N1664265 VSENSE MID N1663951 N1664165 CLAMP_AMP_HI_INA849_OUTAMP
+  PARAMS:  G=500
X_U18           N1663947 N1664179 CLAMP MID GR_SRC_INA849_OUTAMP PARAMS:  GAIN=1 IPOS=70
+  INEG=-70
X_U19           N2052331 N1394706 VOS_DRIFT_INA849_OUTAMP PARAMS:  DC=5U POL=1 DRIFT=1U
X_U20           OUP_OUT VCC VEE ESD_OUT_INA849_OUTAMP
X_U23           N1939580 MID MID N1940296 ZO_SRC_INA849_OUTAMP PARAMS:  GAIN=20 IPOS=35E3
+  INEG=-35E3
X_U4            N995776 N953203 MID N261787 AOL_1_INA849_OUTAMP PARAMS:  GAIN=1E-4 IPOS=.5
+  INEG=-.5
X_U5            N261787 MID MID CLAMP AOL_2_INA849_OUTAMP PARAMS:  GAIN=6.128 IPOS=31.7
+  INEG=-31.7
X_U_OUTAMP_IQN  MID VIMON VEE MID IQ_SRC_INA849_OUTAMP PARAMS:  GAIN=1E-3
X_U_OUTAMP_IQP  VIMON MID MID VCC IQ_SRC_INA849_OUTAMP PARAMS:  GAIN=1E-3
.MODEL R_NOISELESS RES (T_ABS=-273.15)
.ENDS  INA849_OUTAMP
*
.SUBCKT AOL_1_INA849_OUTAMP VC+ VC- IOUT+ IOUT- PARAMS: GAIN=1E-4 IPOS=.5 INEG=-.5
G1 IOUT+ IOUT- VALUE={LIMIT(GAIN*V(VC+,VC-),INEG,IPOS)}
.ENDS  AOL_1_INA849_OUTAMP
*
.SUBCKT AOL_2_INA849_OUTAMP VC+ VC- IOUT+ IOUT- PARAMS: GAIN=20.36E-3 IPOS=0.163 INEG=-0.163
G1 IOUT+ IOUT- VALUE={LIMIT(GAIN*V(VC+,VC-),INEG,IPOS)}
.ENDS  AOL_2_INA849_OUTAMP
*
.SUBCKT CLAMP_AMP_HI_INA849_OUTAMP VC+ VC- VIN COM VO+ VO- PARAMS: G=10
GVO+ COM VO+ VALUE = {IF(V(VIN,COM)>V(VC+,COM),((V(VIN,COM)-V(VC+,COM))*G),0)}
GVO- COM VO- VALUE = {IF(V(VIN,COM)<V(VC-,COM),((V(VC-,COM)-V(VIN,COM))*G),0)}
.ENDS  CLAMP_AMP_HI_INA849_OUTAMP
*
.SUBCKT CLAMP_AMP_LO_INA849_OUTAMP VC+ VC- VIN COM VO+ VO- PARAMS: G=1
GVO+ COM VO+ VALUE = {IF(V(VIN,COM)>V(VC+,COM),((V(VIN,COM)-V(VC+,COM))*G),0)}
GVO- COM VO- VALUE = {IF(V(VIN,COM)<V(VC-,COM),((V(VC-,COM)-V(VIN,COM))*G),0)}
.ENDS  CLAMP_AMP_LO_INA849_OUTAMP
*
.SUBCKT CLAWN_INA849_OUTAMP VC+ VC- IOUT+ IOUT-
G1 IOUT+ IOUT- TABLE {(V(VC+,VC-))} =
+(0, 4.91E-5)
+(4, 1.09E-4)
+(10, 1.66E-4)
+(14, 2.27E-4)
+(18, 3.20E-4)
+(20, 4.56E-4)
+(21, 6.63E-4)
+(22, 9.86E-4)
+(23, 1.42E-3)
+(34, 1.45E-2)
.ENDS  CLAWN_INA849_OUTAMP
*
.SUBCKT CLAWP_INA849_OUTAMP VC+ VC- IOUT+ IOUT-
G1 IOUT+ IOUT- TABLE {(V(VC+,VC-))} =
+(0, 9.41E-5)
+(4, 1.66E-4)
+(10, 2.42E-4)
+(14, 3.41E-4)
+(18, 4.78E-4)
+(20, 5.60E-4)
+(22, 6.72E-4)
+(23, 7.69E-4)
+(24, 9.16E-4)
+(25, 1.11E-3)
+(34, 1.45E-2)
.ENDS  CLAWP_INA849_OUTAMP
*
.SUBCKT CLAW_SRC_INA849_OUTAMP VC+ VC- IOUT+ IOUT- PARAMS: GAIN=1 IPOS=0.226E1 INEG=-0.226E1
G1 IOUT+ IOUT- VALUE={LIMIT(GAIN*V(VC+,VC-),INEG,IPOS)}
.ENDS  CLAW_SRC_INA849_OUTAMP
*
.SUBCKT CL_SRC_INA849_OUTAMP VC+ VC- IOUT+ IOUT- PARAMS: GAIN=1 IPOS=0.452E1 INEG=-0.452E1
G1 IOUT+ IOUT- VALUE={LIMIT(GAIN*V(VC+,VC-),INEG,IPOS)}
.ENDS  CL_SRC_INA849_OUTAMP
*
.SUBCKT ESD_OUT_INA849_OUTAMP OUT VCC VEE
.MODEL ESD_SW VSWITCH(RON=50 ROFF=1E12 VON=500E-3 VOFF=100E-3)
S1 VCC OUT OUT VCC ESD_SW
S2 OUT VEE VEE OUT ESD_SW
.ENDS  ESD_OUT_INA849_OUTAMP
*
.SUBCKT GR_SRC_INA849_OUTAMP VC+ VC- IOUT+ IOUT- PARAMS: GAIN=1 IPOS=0.326E1 INEG=-0.326E1
G1 IOUT+ IOUT- VALUE={LIMIT(GAIN*V(VC+,VC-),INEG,IPOS)}
.ENDS  GR_SRC_INA849_OUTAMP
*
.SUBCKT IQ_SRC_INA849_OUTAMP VC+ VC- IOUT+ IOUT- PARAMS: GAIN=1E-3
G1 IOUT+ IOUT- VALUE={IF( (V(VC+,VC-)<=0),0,GAIN*V(VC+,VC-) )}
.ENDS  IQ_SRC_INA849_OUTAMP
*
.SUBCKT OUTAMP_BLOCK_DC_H_IMON_INA849_OUTAMP 1 2 3 4
H_H_IMON         3 4 VH_H_IMON 1K
VH_H_IMON         1 2 0V
.ENDS  OUTAMP_BLOCK_DC_H_IMON_INA849_OUTAMP
*
.SUBCKT VCM_CLAMP_INA849_OUTAMP VIN+ VIN- IOUT- IOUT+ VP+ VP- PARAMS: GAIN=1
G1 IOUT+ IOUT- VALUE={LIMIT(GAIN*V(VIN+,VIN-),V(VP-,VIN-), V(VP+,VIN-))}
.ENDS  VCM_CLAMP_INA849_OUTAMP
*
.SUBCKT VNSE1_INA849_OUTAMP 1 2 PARAMS: FLW=1 NLF=120 NVR=18
.PARAM GLF={PWR(FLW,0.25)*NLF/1164}
.PARAM RNV={1.184*PWR(NVR,2)}
.MODEL DVN D KF={PWR(FLW,0.5)/1E11} IS=1.0E-16
I1 0 7 10E-3
I2 0 8 10E-3
D1 7 0 DVN
D2 8 0 DVN
E1 3 6 7 8 {GLF}
R1 3 0 1E9
R2 3 0 1E9
R3 3 6 1E9
E2 6 4 5 0 10
R4 5 0 {RNV}
R5 5 0 {RNV}
R6 3 4 1E9
R7 4 0 1E9
E3 1 2 3 4 1
.ENDS  VNSE1_INA849_OUTAMP
*
.SUBCKT VOS_DRIFT_INA849_OUTAMP VOS+ VOS- PARAMS: DC=496.4E-6 POL=1 DRIFT=2E-06
E1 VOS+ VOS- VALUE={DC+POL*DRIFT*(TEMP-27)}
.ENDS  VOS_DRIFT_INA849_OUTAMP
*
.SUBCKT ZO_SRC_INA849_OUTAMP VC+ VC- IOUT+ IOUT- PARAMS: GAIN=200 IPOS=14.5E5 INEG=-14.5E5
G1 IOUT+ IOUT- VALUE={LIMIT(GAIN*V(VC+,VC-),INEG,IPOS)}
.ENDS  ZO_SRC_INA849_OUTAMP
*$
*
*****************************************************************************
.SUBCKT INA849_INAMP INP_IN+ INP_IN- MID VCC VEE INP_OUT
*****************************************************************************
C_C10          N256245 N256255  787.9N
C_C11          MID N257223  43.6P
C_C21          N256265 N256273  3.577P
C_C22          MID N257277  83F
C_C25          CLAMP1 MID  8.204N
C_C28          MID N957967  83F
C_C_VIMON11    VIMON1 MID  1P
G_G12          VSENSE1 MID CLAMP1 MID -1M
G_G15          N256245 MID VSENSE1 N256819 -89
G_G16          N256555 MID N256255 MID -3.505
G_G17          N256265 MID N256573 MID -1
G_G26          N256623 MID N256273 MID -1.022
G_G27          N256659 MID N256643 MID -1
G_G55          N256703 MID N957915 MID -1
R_R136         MID VSENSE1 R_NOISELESS 1K
R_R143         N957915 N256659 R_NOISELESS 9.8K
R_R144         N957967 N957915 R_NOISELESS 10K
R_R34          N256255 N256245 R_NOISELESS 10K
R_R35          MID N256245 R_NOISELESS 1
R_R36          MID N256255 R_NOISELESS 3.992K
R_R38          N256573 N256555 R_NOISELESS 224.1
R_R39          N257223 N256573 R_NOISELESS 10K
R_R41          MID N256265 R_NOISELESS 1
R_R46          MID N256555 R_NOISELESS 1
R_R67          N256273 N256265 R_NOISELESS 10K
R_R68          MID N256623 R_NOISELESS 1
R_R69          MID N256273 R_NOISELESS 445K
R_R70          N256643 N256623 R_NOISELESS 9.8K
R_R71          N257277 N256643 R_NOISELESS 10K
R_R72          MID N256659 R_NOISELESS 1
R_R75          MID N256703 R_NOISELESS 1
R_R78          MID N261786 R_NOISELESS 1MEG
R_R79          MID CLAMP1 R_NOISELESS 1MEG
R_RDUMMY1      MID N256819 R_NOISELESS 575
R_RIN1         N928127 INP_IN+ R_NOISELESS 10M
R_RIN2         N928131 INP_IN- R_NOISELESS 10M
R_RX1          N256819 N256703 R_NOISELESS 5.75K
R_R_VIMON11    N970369 VIMON1 R_NOISELESS 100
R_R_VIMON12    MID N970369 R_NOISELESS 1T
X_H_IMON11     N256819 INP_OUT N970369 MID INA849_INAMP_H_IMON11
X_U2           N928127 N928131 MID N261786 AOL_1_INA849_INAMP PARAMS:  GAIN=1E-4 IPOS=.5
+  INEG=-.5
X_U3           N261786 MID MID CLAMP1 AOL_2_INA849_INAMP PARAMS:  GAIN=8.848E-3 IPOS=4 INEG=-4
X_U_INAMP_IQN  MID VIMON1 VEE MID IQ_SRC_INA849_INAMP PARAMS:  GAIN=1E-3
X_U_INAMP_IQP  VIMON1 MID MID VCC IQ_SRC_INA849_INAMP PARAMS:  GAIN=1E-3
.MODEL R_NOISELESS RES (T_ABS=-273.15)
.ENDS  INA849_INAMP
*
.SUBCKT AOL_1_INA849_INAMP VC+ VC- IOUT+ IOUT- PARAMS: GAIN=1E-4 IPOS=.5 INEG=-.5
G1 IOUT+ IOUT- VALUE={LIMIT(GAIN*V(VC+,VC-),INEG,IPOS)}
.ENDS  AOL_1_INA849_INAMP
*
.SUBCKT AOL_2_INA849_INAMP VC+ VC- IOUT+ IOUT- PARAMS: GAIN=20.36E-3 IPOS=0.163 INEG=-0.163
G1 IOUT+ IOUT- VALUE={LIMIT(GAIN*V(VC+,VC-),INEG,IPOS)}
.ENDS  AOL_2_INA849_INAMP
*
.SUBCKT INA849_INAMP_H_IMON11 1 2 3 4
H_H_IMON11         3 4 VH_H_IMON11 1K
VH_H_IMON11         1 2 0V
.ENDS  INA849_INAMP_H_IMON11
*
.SUBCKT IQ_SRC_INA849_INAMP VC+ VC- IOUT+ IOUT- PARAMS: GAIN=1E-3
G1 IOUT+ IOUT- VALUE={IF( (V(VC+,VC-)<=0),0,GAIN*V(VC+,VC-) )}
.ENDS  IQ_SRC_INA849_INAMP
*
