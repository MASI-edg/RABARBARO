*$
* OPA161x
*****************************************************************************
* (C) Copyright 2022 Texas Instruments Incorporated. All rights reserved.                                            
*****************************************************************************
** This model is designed as an aid for customers of Texas Instruments.
** TI and its licensors and suppliers make no warranties, either expressed
** or implied, with respect to this model, including the warranties of 
** merchantability or fitness for a particular purpose.  The model is
** provided solely on an "as is" basis.  The entire risk as to its quality
** and performance is with the customer
*****************************************************************************
*
* This model is subject to change without notice. Texas Instruments
* Incorporated is not responsible for updating this model.
*
*****************************************************************************
*
** Released by: Online Design Tools, Texas Instruments Inc.
* Part: OPA161x
* Date: 24AUG2022
* Model Type: Generic (suitable for all analysis types)
* EVM Order Number: N/A 
* EVM Users Guide:  N/A 
* Datasheet: SBOS450C -JULY 2009-REVISED AUGUST 2014 
* Created with Green-Williams-Lis Op Amp Macro-model Architecture
*
* Model Version: Final 1.5
*
*****************************************************************************
*
* Updates:
*
* Final 1.5
* 1. Moved R_NOISELESS .model inside OPA161x subckt.
* 2. Updated PSpice Symbol.
*
* Final 1.4
* 1. Updated the current direction(i.e. IOUT- IOUT+) of IQ_SRC block to 
*    resolve Iout current direction issue.
* 2. Added R_DIFF element in the model.
*
* Final 1.3
* 1. Modified the capacitor(C14) value from 1F to 2.5uF in GND Float-IQ block  
*    to resolve the convergence issue in single and asymmetric supply test.
* 2. Remodeled CMRR last stage to resolve the issue in Voltage Noise result
*    while simulating in PSpice.
* 3. Updated the model name from OPA1611 to OPA161x.
*
* Final 1.2
* 1. VOS drift feature is added 
* 2. Added Unique subckt name, removed Claw ABS.
*
* Final 1.1 
* Release to Web.
*
*****************************************************************************
* Model Usage Notes:
* 1. The following parameters are modeled: 
*    a. OPEN-LOOP GAIN AND PHASE VS. FREQUENCY  WITH RL, CL EFFECTS (Aol)
*    b. UNITY GAIN BANDWIDTH (GBW)
*    c. INPUT COMMON-MODE REJECTION RATIO VS. FREQUENCY (CMRR)
*    d. POWER SUPPLY REJECTION RATIO VS. FREQUENCY (PSRR)
*    e. DIFFERENTIAL INPUT IMPEDANCE (Zid)
*    f. COMMON-MODE INPUT IMPEDANCE (Zic)
*    g. OPEN-LOOP OUTPUT IMPEDANCE VS. FREQUENCY (Zo)
*    h. OUTPUT CURRENT THROUGH THE SUPPLY (Iout)
*    i. INPUT VOLTAGE NOISE DENSITY VS. FREQUENCY (en)
*    j. INPUT CURRENT NOISE DENSITY VS. FREQUENCY (in)
*    k. OUTPUT VOLTAGE SWING vs. OUTPUT CURRENT (Vo)
*    l. SHORT-CIRCUIT OUTPUT CURRENT (Isc)
*    m. QUIESCENT CURRENT (Iq)
*    n. SETTLING TIME VS. CAPACITIVE LOAD (ts)
*    o. SLEW RATE (SR)
*    p. SMALL SIGNAL OVERSHOOT VS. CAPACITIVE LOAD
*    q. LARGE SIGNAL RESPONSE
*    r. OVERLOAD RECOVERY TIME (tor)
*    s. INPUT BIAS CURRENT (Ib)
*    t. INPUT OFFSET CURRENT (Ios)
*    u. INPUT OFFSET VOLTAGE (Vos)
*    v. INPUT OFFSET VOLTAGE VS. TEMPERATURE (Vos Drift)
*    w. INPUT COMMON-MODE VOLTAGE RANGE (Vcm)
*    x. INPUT OFFSET VOLTAGE VS. INPUT COMMON-MODE VOLTAGE (Vos vs. Vcm)
*    y. INPUT/OUTPUT ESD CELLS (ESDin, ESDout)
* 2. OPA161x model is available in single core(OPA1611) and dual 
*    core(OPA1612).
*****************************************************************************
.SUBCKT OPA161x IN+ IN- VCC VEE OUT  
*****************************************************************************
C_C1          N24458 N24659  22.044F 
C_C10         N37029 N37037  117.6646N 
C_C11         MID N39473  1.175576P 
C_C12         N39884 N39892  413.8029F 
C_C13         0 N2392253  1F 
C_C14         0 N2392113  2.5U 
C_C15         0 N2392293  1F 
C_C16         MID N56849  1F 
C_C17         MID N57325  1F 
C_C18         MID N59747  1F 
C_C19         MID N59865  1F 
C_C2          N25921 N25929  214.32P 
C_C20         MID N65579  1F 
C_C21         MID N65697  1F 
C_C22         MID N68774  1F 
C_C23         N72398 MID  1F 
C_C24         MID N72391  1F 
C_C25         MID N81574  1P 
C_C26         MID N81664  1P 
C_C27         MID SW_OL_OPA161x  1N 
C_C28         VCLP MID  1P 
C_C29         VIMON MID  1P 
C_C3          N27785 N27793  318.31P 
C_C30         VOUT_S MID  1P 
C_C31         N2402147 N2402155  220.4P 
C_C32         MID N2419074  23.15998F 
C_C33         N2423000 N36262  1.428314P 
C_C4          N32347 MID  1F 
C_C5          CLAMP MID  925.2513P 
C_C6          N34005 N34013  106.1033F 
C_C_COM0      ESDP MID  2P 
C_C_COM1      MID ESDN  2P 
C_C_DIFF      ESDN ESDP  8P 
E_E1          MID 0 N2392113 0 1
E_E2          N158495 MID CL_CLAMP MID 1
E_E3          N161937 MID OUT MID 1
G_G1          N24458 MID ESDP MID -162.65U
G_G12         CLAW_CLAMP MID N36262 MID -1M
G_G13         CL_CLAMP MID CLAW_CLAMP MID -1M
G_G15         N37029 MID CL_CLAMP N45999 -89.0524
G_G16         N39124 MID N37037 MID -270.7824
G_G17         N39884 MID N39417 MID -1
G_G18         VCC_B 0 VCC 0 -1
G_G19         VEE_B 0 VEE 0 -1
G_G2          N25415 N25397 N25248 MID -1M
G_G20         VCC_CLP MID N72398 MID -1M
G_G21         VEE_CLP MID N72391 MID -1M
G_G22         N1356345 MID N1356333 MID -1
G_G23         N1356409 MID N1356429 MID -1
G_G24         N2402147 MID N24659 MID -1
G_G25         N25248 MID N2402155 MID -140.5
G_G26         N2419074 MID VSENSE MID -1U
G_G27         N2423000 MID N34013 MID -21.5263
G_G3          N25921 MID VEE_B MID -115.72M
G_G4          N27785 MID VCC_B MID -121.95M
G_G5          N28678 N28438 N27793 N25929 -1M
G_G6          VSENSE MID CLAMP MID -1M
G_G8          N34005 MID N2419074 MID -21.5263
I_I_B         N24207 MID DC 60N  
I_I_OS        ESDN MID DC 35N  
I_I_Q         VCC VEE DC 3.6M  
R_R1          IN+ ESDP R_NOISELESS 10M
R_R10         MID N25921 R_NOISELESS 1
R_R11         MID N25929 R_NOISELESS 79.383
R_R12         N27793 N27785 R_NOISELESS 100MEG
R_R13         MID N27785 R_NOISELESS 1
R_R14         MID N27793 R_NOISELESS 74.0813
R_R15         N28438 N25415 R_NOISELESS 1M
R_R16         N28678 N28438 R_NOISELESS 1K
R_R17         N31303 ESDN R_NOISELESS 1M
R_R18         MID N31389 R_NOISELESS 1T
R_R19         MID N31737 R_NOISELESS 1T
R_R2          IN- ESDN R_NOISELESS 10M
R_R20         N32236 MID R_NOISELESS 1
R_R21         N32347 N32236 R_NOISELESS 1M
R_R22         MID N32510 R_NOISELESS 1MEG
R_R23         MID CLAMP R_NOISELESS 1MEG
R_R24         MID VSENSE R_NOISELESS 1K
R_R25         N34013 N34005 R_NOISELESS 10K
R_R26         MID N34005 R_NOISELESS 1
R_R27         MID N34013 R_NOISELESS 487.1795
R_R3          ESDP MID R_NOISELESS 1T
R_R32         MID CLAW_CLAMP R_NOISELESS 1K
R_R33         MID CL_CLAMP R_NOISELESS 1K
R_R34         N37037 N37029 R_NOISELESS 10K
R_R35         MID N37029 R_NOISELESS 1
R_R36         MID N37037 R_NOISELESS 37.0669
R_R37         MID N39124 R_NOISELESS 1
R_R38         N39417 N39124 R_NOISELESS 1.312633MEG
R_R39         N39473 N39417 R_NOISELESS 10K
R_R4          MID ESDN R_NOISELESS 1T
R_R40         N39892 N39884 R_NOISELESS 10K
R_R41         MID N39884 R_NOISELESS 1
R_R42         MID N39892 R_NOISELESS 9.268057
R_R43         MID N46041 R_NOISELESS 1
R_R46         VCC_B 0 R_NOISELESS 1
R_R47         VCC_B N2392253 R_NOISELESS 1M
R_R48         N2392253 N2392113 R_NOISELESS 1MEG
R_R49         N2392113 0 R_NOISELESS 1T
R_R5          MID N24458 R_NOISELESS 1
R_R50         N2392113 N2392293 R_NOISELESS 1MEG
R_R51         N2392293 VEE_B R_NOISELESS 1M
R_R52         VEE_B 0 R_NOISELESS 1
R_R53         VCC_CLP MID R_NOISELESS 1T
R_R54         N55560 MID R_NOISELESS 1
R_R55         N56849 N55560 R_NOISELESS 1M
R_R56         VEE_CLP MID R_NOISELESS 1T
R_R57         N57321 MID R_NOISELESS 1
R_R58         N57325 N57321 R_NOISELESS 1M
R_R59         N59739 MID R_NOISELESS 1T
R_R6          N24659 N24458 R_NOISELESS 100MEG
R_R60         N59743 MID R_NOISELESS 1
R_R61         N59747 N59743 R_NOISELESS 1M
R_R62         N59865 N59881 R_NOISELESS 1M
R_R63         N59905 MID R_NOISELESS 1T
R_R64         N59881 MID R_NOISELESS 1
R_R65         N65567 MID R_NOISELESS 1T
R_R66         N65575 MID R_NOISELESS 1
R_R67         N65579 N65575 R_NOISELESS 1M
R_R68         N65697 N65713 R_NOISELESS 1M
R_R69         N65737 MID R_NOISELESS 1T
R_R7          MID N24659 R_NOISELESS 716.778969K
R_R70         N65713 MID R_NOISELESS 1
R_R71         N68774 VSENSE R_NOISELESS 1M
R_R72         VCC_B N72064 R_NOISELESS 1K
R_R73         N72064 N72398 R_NOISELESS 1M
R_R74         N72073 VEE_B R_NOISELESS 1K
R_R75         N72073 N72391 R_NOISELESS 1M
R_R76         MID VCC_CLP R_NOISELESS 1K
R_R77         VEE_CLP MID R_NOISELESS 1K
R_R78         N1356409 MID R_NOISELESS 1
R_R79         N1356345 MID R_NOISELESS 1
R_R8          N25415 N25397 R_NOISELESS 1K
R_R80         V11 N81574 R_NOISELESS 100
R_R81         V12 N81664 R_NOISELESS 100
R_R82         N81756 MID R_NOISELESS 1
R_R83         N81756 SW_OL_OPA161x R_NOISELESS 100
R_R84         N158495 VCLP R_NOISELESS 100
R_R85         N2402155 N2402147 R_NOISELESS 10K
R_R86         MID N2402147 R_NOISELESS 1
R_R87         MID N2402155 R_NOISELESS 71.69
R_R88         MID N25248 R_NOISELESS 1
R_R89         MID N2419074 R_NOISELESS 1MEG
R_R9          N25929 N25921 R_NOISELESS 100MEG
R_R90         N36262 N2423000 R_NOISELESS 10K
R_R91         MID N2423000 R_NOISELESS 1
R_R92         MID N36262 R_NOISELESS 487.1795
R_RDUMMY      MID N45999 R_NOISELESS 1.41K
R_R_DIFF      ESDN ESDP R_NOISELESS 100MEG
R_RX          N45999 N46041 R_NOISELESS 14.1K
R_RX1         MID N161737 R_NOISELESS 1T
R_RX2         VIMON N161737 R_NOISELESS 100
R_RX3         MID N161937 R_NOISELESS 1T
R_RX4         VOUT_S N161937 R_NOISELESS 100
V_VCM_MAX     N31389 VCC_B -2
V_VCM_MIN     N31737 VEE_B 2
V_V_GRN       N65737 MID -47
V_V_GRP       N65567 MID 48
V_V_ISCN      N59905 MID -47
V_V_ISCP      N59739 MID 49.8
V_V_ORN       N1356333 VCLP -13.759
V_V_ORP       N1356429 VCLP 13.6794
X_H1          N45999 OUT N161737 MID BLOCK_DC_H1_OPA161x 
X_H2          N1356115 N1356409 V12 MID BLOCK_DC_H2_OPA161x 
X_H3          N1356061 N1356345 V11 MID BLOCK_DC_H3_OPA161x 
X_S1          N1356061 CLAMP N1356061 CLAMP BLOCK_DC_S1_OPA161x 
X_S2          CLAMP N1356115 CLAMP N1356115 BLOCK_DC_S2_OPA161x 
X_U1          ESDP N24207 VNSE_OPA161x PARAMS: FLW=0.1 GLF=0.01152 RNV=1.8205
X_U10         VCC_CLP VEE_CLP VOUT_S MID N55560 N57321 CLAMP_AMP_LO_OPA161x PARAMS: G=1
X_U11         N59739 N59905 VIMON MID N59743 N59881 CLAMP_AMP_LO_OPA161x PARAMS: G=1
X_U12         N65567 N65737 N68774 MID N65575 N65713 CLAMP_AMP_HI_OPA161x PARAMS: G=10
X_U16         MID N81756 N81574 N81664 OL_SENSE_OPA161x
X_U18         VIMON MID N72064 VCC_B CLAWP_OPA161x
X_U19         MID VIMON VEE_B N72073 CLAWN_OPA161x
X_U20         ESDN ESDP ESD_BB_OPA161x
X_U21         OUT VCC VEE ESD_OUT_OPA161x
X_U22         N59747 N59865 CL_CLAMP MID CL_SRC_OPA161x PARAMS: GAIN=1 IPOS=0.2016E1
+  INEG=-0.1974E1
X_U23         N65579 N65697 CLAMP MID GR_SRC_OPA161x PARAMS: GAIN=1 IPOS=0.056064E1
+  INEG=-0.056064E1
X_U25         SW_OL_OPA161x MID N37029 N37037 SW_OL_OPA161x PARAMS:
X_U26         VIMON MID MID VCC IQ_SRC_OPA161x PARAMS: GAIN=1E-3
X_U27         MID VIMON VEE MID IQ_SRC_OPA161x PARAMS: GAIN=1E-3
X_U30         N32347 N31303 MID N32510 AOL_1_OPA161x PARAMS: GAIN=1E-4 IPOS=.5 INEG=-.5
X_U31         N32510 MID MID CLAMP AOL_2_OPA161x PARAMS: GAIN=0.0053649 IPOS=0.025232
+  INEG=-0.025211
X_U32         N39892 MID MID N46041 ZO_SRC_OPA161x PARAMS: GAIN=1079.9748 IPOS=1551E4
+  INEG=-1748.4E4
X_U35         N56849 N57325 CLAW_CLAMP MID CLAW_SRC_OPA161x PARAMS: GAIN=1
+  IPOS=0.1008E1 INEG=-0.0987E1
X_U36         N24207 MID FEMT_OPA161x PARAMS: FLWF=0.1 GLFF=19.0969 RNVF=3.366E6
X_U37         ESDN MID FEMT_OPA161x PARAMS: FLWF=0.1 GLFF=19.0969 RNVF=3.366E6
X_U4          N25397 N24207 VOS_DRIFT_OPA161x PARAMS: DC=9.729E-05 POL=1 DRIFT=1E-06
X_U5          ESDN ESDP VCC VEE ESD_IN_OPA161x
X_U6          N28678 MID N32236 MID N31389 N31737 VCM_CLAMP_OPA161x PARAMS: GAIN=1
.MODEL R_NOISELESS RES (T_ABS=-273.15)
.ENDS OPA161x
*
.SUBCKT BLOCK_DC_H1_OPA161x 1 2 3 4  
H_H1         3 4 VH_H1 1K
VH_H1         1 2 0V
.ENDS  BLOCK_DC_H1_OPA161x
*
.SUBCKT BLOCK_DC_H2_OPA161x 1 2 3 4  
H_H2         3 4 VH_H2 1
VH_H2         1 2 0V
.ENDS  BLOCK_DC_H2_OPA161x
*
.SUBCKT BLOCK_DC_H3_OPA161x 1 2 3 4  
H_H3         3 4 VH_H3 -1
VH_H3         1 2 0V
.ENDS  BLOCK_DC_H3_OPA161x
*
.SUBCKT BLOCK_DC_S1_OPA161x 1 2 3 4  
S_S1         3 4 1 2 _S1
RS_S1         1 2 1G
.MODEL         _S1 VSWITCH ROFF=1E12 RON=10M VOFF=0.0V VON=10MV
.ENDS  BLOCK_DC_S1_OPA161x
*
.SUBCKT BLOCK_DC_S2_OPA161x 1 2 3 4  
S_S2         3 4 1 2 _S2
RS_S2         1 2 1G
.MODEL         _S2 VSWITCH ROFF=1E12 RON=10M VOFF=0.0V VON=10MV
.ENDS  BLOCK_DC_S2_OPA161x
*
.SUBCKT AOL_1_OPA161x VC+ VC- IOUT+ IOUT- PARAMS: GAIN=1E-4 IPOS=.5 INEG=-.5
G1 IOUT+ IOUT- VALUE={LIMIT(GAIN*V(VC+,VC-),INEG,IPOS)}
.ENDS  AOL_1_OPA161x
*
.SUBCKT AOL_2_OPA161x VC+ VC- IOUT+ IOUT- PARAMS: GAIN=0.0053649 IPOS=0.025232 INEG=-0.025211
G1 IOUT+ IOUT- VALUE={LIMIT(GAIN*V(VC+,VC-),INEG,IPOS)}
.ENDS  AOL_2_OPA161x
*
.SUBCKT CLAMP_AMP_HI_OPA161x VC+ VC- VIN COM VO+ VO- PARAMS: G=10
GVO+ COM VO+ VALUE = {IF(V(VIN,COM)>V(VC+,COM),((V(VIN,COM)-V(VC+,COM))*G),0)}
GVO- COM VO- VALUE = {IF(V(VIN,COM)<V(VC-,COM),((V(VC-,COM)-V(VIN,COM))*G),0)}
.ENDS  CLAMP_AMP_HI_OPA161x
*
.SUBCKT CLAMP_AMP_LO_OPA161x VC+ VC- VIN COM VO+ VO- PARAMS: G=1
GVO+ COM VO+ VALUE = {IF(V(VIN,COM)>V(VC+,COM),((V(VIN,COM)-V(VC+,COM))*G),0)}
GVO- COM VO- VALUE = {IF(V(VIN,COM)<V(VC-,COM),((V(VC-,COM)-V(VIN,COM))*G),0)}
.ENDS  CLAMP_AMP_LO_OPA161x
*
.SUBCKT CLAWN_OPA161x VC+ VC- IOUT+ IOUT-
G1 IOUT+ IOUT- TABLE {(V(VC+,VC-))} =
+(0, 2.1349E-4)
+(45.4769, 0.0008314)
+(46.5224, 0.00085953)
+(47, 0.0010745)
.ENDS  CLAWN_OPA161x
*
.SUBCKT CLAWP_OPA161x VC+ VC- IOUT+ IOUT-
G1 IOUT+ IOUT- TABLE {(V(VC+,VC-))} =
+(0, 2.1334E-4)
+(48.1473, 0.001)
+(49.2541, 0.0012)
+(49.8, 0.0013)
.ENDS  CLAWP_OPA161x
*
.SUBCKT CLAW_SRC_OPA161x VC+ VC- IOUT+ IOUT- PARAMS: GAIN=1 IPOS=0.1008E1 INEG=-0.0987E1
G1 IOUT+ IOUT- VALUE={LIMIT(GAIN*V(VC+,VC-),INEG,IPOS)}
.ENDS  CLAW_SRC_OPA161x
*
.SUBCKT CL_SRC_OPA161x VC+ VC- IOUT+ IOUT- PARAMS: GAIN=1 IPOS=0.2016E1 INEG=-0.1974E1
G1 IOUT+ IOUT- VALUE={LIMIT(GAIN*V(VC+,VC-),INEG,IPOS)}
.ENDS  CL_SRC_OPA161x
*
.SUBCKT ESD_BB_OPA161x ESDN ESDP
.MODEL ESD_SW VSWITCH(RON=50 ROFF=1E12 VON=700E-3 VOFF=0)
S1 ESDN ESDP ESDN ESDP ESD_SW
S2 ESDP ESDN ESDP ESDN ESD_SW
.ENDS  ESD_BB_OPA161x
*
.SUBCKT ESD_IN_OPA161x ESDN ESDP VCC VEE
.MODEL ESD_SW VSWITCH(RON=50 ROFF=1E12 VON=500E-3 VOFF=100E-3)
S1 ESDN VCC ESDN VCC ESD_SW
S2 ESDP VCC ESDP VCC ESD_SW
S3 VEE ESDN VEE ESDN ESD_SW
S4 VEE ESDP VEE ESDP ESD_SW
.ENDS  ESD_IN_OPA161x
*
.SUBCKT ESD_OUT_OPA161x OUT VCC VEE
.MODEL ESD_SW VSWITCH(RON=50 ROFF=1E12 VON=500E-3 VOFF=100E-3)
S1 OUT VCC OUT VCC ESD_SW
S2 VEE OUT VEE OUT ESD_SW
.ENDS  ESD_OUT_OPA161x
*
.SUBCKT FEMT_OPA161x 1 2 PARAMS: FLWF=0.1 GLFF=19.0969 RNVF=3.366E6
.MODEL DVNF D KF={PWR(FLWF,0.5)/1E11} IS=1.0E-16
I1 0 7 10E-3
I2 0 8 10E-3
D1 7 0 DVNF
D2 8 0 DVNF
E1 3 6 7 8 {GLFF}
R1 3 0 1E9
R2 3 0 1E9
R3 3 6 1E9
E2 6 4 5 0 10
R4 5 0 {RNVF}
R5 5 0 {RNVF}
R6 3 4 1E9
R7 4 0 1E9
G1 1 2 3 4 1E-6
.ENDS  FEMT_OPA161x
*
.SUBCKT GR_SRC_OPA161x VC+ VC- IOUT+ IOUT- PARAMS: GAIN=1 IPOS=0.056064E1 INEG=-0.056064E1
G1 IOUT+ IOUT- VALUE={LIMIT(GAIN*V(VC+,VC-),INEG,IPOS)}
.ENDS  GR_SRC_OPA161x
*
.SUBCKT IQ_SRC_OPA161x VC+ VC- IOUT+ IOUT- PARAMS: GAIN=1E-3
G1 IOUT- IOUT+ VALUE={IF( (V(VC+,VC-)<=0),0,GAIN*V(VC+,VC-) )}
.ENDS  IQ_SRC_OPA161x
*
.SUBCKT OL_SENSE_OPA161x COM SW+ OLN OLP
GSW+ COM SW+ VALUE = {IF((V(OLN,COM)>10E-3 | V(OLP,COM)>10E-3),1,0)}
.ENDS  OL_SENSE_OPA161x
*
.SUBCKT SW_OL_OPA161x SW_OL_OPA161x MID CAP_L CAP_R
.MODEL OL_SW VSWITCH(RON=1E-3 ROFF=1E12 VON=900E-3 VOFF=800E-3)
S1 CAP_L CAP_R SW_OL_OPA161x MID OL_SW
.ENDS  SW_OL_OPA161x
*
.SUBCKT VCM_CLAMP_OPA161x VIN+ VIN- IOUT- IOUT+ VP+ VP- PARAMS: GAIN=1
G1 IOUT+ IOUT- VALUE={LIMIT(GAIN*V(VIN+,VIN-),V(VP-,VIN-), V(VP+,VIN-))}
.ENDS  VCM_CLAMP_OPA161x
*
.SUBCKT VNSE_OPA161x 1 2 PARAMS: FLW=0.1 GLF=0.01152 RNV=1.8205
.MODEL DVN D KF={PWR(FLW,0.5)/1E11} IS=1.0E-16
I1 0 7 10E-3
I2 0 8 10E-3
D1 7 0 DVN
D2 8 0 DVN
E1 3 6 7 8 {GLF}
R1 3 0 1E9
R2 3 0 1E9
R3 3 6 1E9
E2 6 4 5 0 10
R4 5 0 {RNV}
R5 5 0 {RNV}
R6 3 4 1E9
R7 4 0 1E9
E3 1 2 3 4 1
.ENDS  VNSE_OPA161x
*
.SUBCKT VOS_DRIFT_OPA161x VOS+ VOS- PARAMS: DC=9.729E-05 POL=1 DRIFT=1E-06
E1 VOS+ VOS- VALUE={DC+POL*DRIFT*(TEMP-27)}
.ENDS  VOS_DRIFT_OPA161x
*
.SUBCKT ZO_SRC_OPA161x VC+ VC- IOUT+ IOUT- PARAMS: GAIN=1079.9748 IPOS=1551E4 INEG=-1748.4E4
G1 IOUT+ IOUT- VALUE={LIMIT(GAIN*V(VC+,VC-),INEG,IPOS)}
.ENDS  ZO_SRC_OPA161x
*
